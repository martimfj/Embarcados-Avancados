// niosHello_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module niosHello_tb (
	);

	wire    nioshello_inst_clk_bfm_clk_clk;       // niosHello_inst_clk_bfm:clk -> [niosHello_inst:clk_clk, niosHello_inst_reset_bfm:clk]
	wire    nioshello_inst_reset_bfm_reset_reset; // niosHello_inst_reset_bfm:reset -> niosHello_inst:reset_reset_n

	niosHello nioshello_inst (
		.clk_clk       (nioshello_inst_clk_bfm_clk_clk),       //   clk.clk
		.keys_export   (),                                     //  keys.export
		.leds_name     (),                                     //  leds.name
		.reset_reset_n (nioshello_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nioshello_inst_clk_bfm (
		.clk (nioshello_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nioshello_inst_reset_bfm (
		.reset (nioshello_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nioshello_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
